module ALU_Control
(
	input [1:0] ALUOp, 
	input [3:0] Funct,
	output reg [3:0] Operation
);

	always @ (ALUOp or Funct)
	begin
		case(ALUOp)
			2'b00: begin
			case(Funct)
			     2'b0001: Operation = 4'b1111;
			     default: Operation = 4'b0010;
			endcase
			end
			2'b01: 
			begin 
			case(Funct)
			    4'b0100:Operation = 4'b1110; //Generating new control signal in case of blt
			    default:Operation = 4'b0110;			    
			endcase
			end
			2'b10:
			begin 
			case(Funct)
				4'b0000: Operation = 4'b0010;
				4'b1000: Operation = 4'b0110;
				4'b0111: Operation = 4'b0000;
				4'b0110: Operation = 4'b0001;
			endcase
			end
		endcase
	end
	
endmodule
